/// INicio